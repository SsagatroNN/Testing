module alu #(
    parameter D_WIDTH = 32
) (
    input logic alusrc,
    input logic [2:0] aluctrl,


endmodule
