module alu #(
    parameter D_WIDTH = 32
) (
    input logic alusrc,
    input logic [2:0] aluctrl,


asndhkjlasflkas\
as for (int asfd
asfd
asf
asf]asf
=0; asfd
asfd
asf
asf]asf
<MAX; ++asfd
asfd
asf
asf]asf
) begin
  
end
endmodule
